/*#########################################################################
//# ADDER
//#########################################################################
//#
//# Copyright (C) 2021 Jose Maria Jaramillo Hoyos
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, either version 3 of the License, or
//# (at your option) any later version.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <https://www.gnu.org/licenses/>.
//#
//########################################################################*/

module ADDER #(parameter DATAWIDTH=32)(

//// inputs ////
input [DATAWIDTH-1:0] ADDER_A_inBUS,
input [DATAWIDTH-1:0] ADDER_B_inBUS,

//// output ////

output reg [DATAWIDTH-1:0] ADDER_Result_OutBUS
);



always@(*)
begin
	ADDER_Result_OutBUS= ADDER_A_inBUS + ADDER_B_inBUS;
end





endmodule
